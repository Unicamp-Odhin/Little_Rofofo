module Little_Rofofo #(
    parameter BOOT_ADDRESS = 32'h00000000,
    parameter DATA_WIDTH   = 32'd32,
    parameter ADDR_WIDTH   = 32'd32,
) (
    input logic clk,
    input logic rst_n
);
    
endmodule
