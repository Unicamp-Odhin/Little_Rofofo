module top (
    input  logic clk,
    input  logic rst_n,

    output logic rx,
    input  logic tx,

    output logic [7:0]led,
    inout  logic [5:0]gpios
);



endmodule
